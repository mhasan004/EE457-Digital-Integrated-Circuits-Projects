*** SPICE deck for cell XOR_2{sch} from library Proj2
*** Created on Tue Mar 17, 2020 00:23:25
*** Last revised on Tue Mar 17, 2020 01:00:52
*** Written on Tue Mar 17, 2020 01:01:53 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: XOR_2{sch}
Mnmos@0 net@38 A net@41 gnd NMOS L=0.35U W=1.75U
Mnmos@1 net@38 net@123 net@47 gnd NMOS L=0.35U W=1.75U
Mnmos@2 net@123 A gnd gnd NMOS L=0.35U W=1.75U
Mnmos@3 net@41 net@95 gnd gnd NMOS L=0.35U W=1.75U
Mnmos@4 net@47 B gnd gnd NMOS L=0.35U W=1.75U
Mnmos@5 net@95 B gnd gnd NMOS L=0.35U W=1.75U
Mnmos@6 out net@38 gnd gnd NMOS L=0.35U W=1.75U
Mpmos@0 net@27 A vdd vdd PMOS L=0.35U W=1.75U
Mpmos@1 net@38 net@123 net@27 vdd PMOS L=0.35U W=1.75U
Mpmos@2 net@123 A vdd vdd PMOS L=0.35U W=3.5U
Mpmos@3 net@27 net@95 vdd vdd PMOS L=0.35U W=1.75U
Mpmos@4 net@38 B net@27 vdd PMOS L=0.35U W=1.75U
Mpmos@5 net@95 B vdd vdd PMOS L=0.35U W=3.5U
Mpmos@6 out net@38 vdd vdd PMOS L=0.35U W=3.5U

* Spice Code nodes in cell cell 'XOR_2{sch}'
VDD VDD 0 DC 3.3
VGND GND 0 DC 0
vin A 0 PULSE(0 3.3 0 1ns 1ns 38ns 80ns)
vin2 B 0 PULSE(0 3.3 0 1ns 1ns 18ns 40ns)
cload out 0 250fF
.tran 0 80n
.include C:\Electric\C5_models.txt
.END

*** SPICE deck for cell NOR_2{sch} from library project_1
*** Created on Tue Mar 03, 2020 18:05:36
*** Last revised on Tue Mar 03, 2020 18:31:41
*** Written on Tue Mar 03, 2020 19:45:12 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: NOR_2{sch}
Mnmos@0 out A gnd gnd NMOS L=0.35U W=1.75U
Mnmos@1 out B gnd gnd NMOS L=0.35U W=1.75U
Mpmos@2 net@58 A vdd vdd PMOS L=0.35U W=1.75U
Mpmos@3 out B net@58 vdd PMOS L=0.35U W=1.75U

* Spice Code nodes in cell cell 'NOR_2{sch}'
VDD VDD 0 DC 3.3
VGND GND 0 DC 0
vin A 0 PULSE(0 3.3 0 1ns 1ns 38ns 80ns)
vin2 B 0 PULSE(0 3.3 0 1ns 1ns 18ns 40ns)
cload out 0 250fF
.tran 0 80n
.include C:\Electric\C5_models.txt
.END

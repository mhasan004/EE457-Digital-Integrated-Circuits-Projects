*** SPICE deck for cell Two_bit_adder2{sch} from library Proj2
*** Created on Tue Mar 17, 2020 22:05:22
*** Last revised on Tue Mar 17, 2020 22:37:50
*** Written on Tue Mar 17, 2020 22:37:54 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Proj2__NAND_2 FROM CELL NAND_2{sch}
.SUBCKT Proj2__NAND_2 A B out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out A net@22 gnd NMOS L=0.35U W=1.75U
Mnmos@1 out A vdd vdd PMOS L=0.35U W=1.75U
Mnmos@2 net@22 B gnd gnd NMOS L=0.35U W=1.75U
Mpmos@1 out B vdd vdd PMOS L=0.35U W=1.75U
.ENDS Proj2__NAND_2

*** SUBCIRCUIT Proj2__XOR_2 FROM CELL XOR_2{sch}
.SUBCKT Proj2__XOR_2 A B out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@38 A net@41 gnd NMOS L=0.35U W=1.75U
Mnmos@1 net@38 net@128 net@47 gnd NMOS L=0.35U W=1.75U
Mnmos@2 net@128 A gnd gnd NMOS L=0.35U W=1.75U
Mnmos@3 net@41 net@113 gnd gnd NMOS L=0.35U W=1.75U
Mnmos@4 net@47 B gnd gnd NMOS L=0.35U W=1.75U
Mnmos@5 net@113 B gnd gnd NMOS L=0.35U W=1.75U
Mnmos@6 out net@38 gnd gnd NMOS L=0.35U W=1.75U
Mpmos@0 net@27 A vdd vdd PMOS L=0.35U W=1.75U
Mpmos@1 net@38 net@128 net@27 vdd PMOS L=0.35U W=1.75U
Mpmos@2 net@128 A vdd vdd PMOS L=0.35U W=3.5U
Mpmos@3 net@27 net@113 vdd vdd PMOS L=0.35U W=1.75U
Mpmos@4 net@38 B net@27 vdd PMOS L=0.35U W=1.75U
Mpmos@5 net@113 B vdd vdd PMOS L=0.35U W=3.5U
Mpmos@6 out net@38 vdd vdd PMOS L=0.35U W=3.5U
.ENDS Proj2__XOR_2

.global gnd vdd

*** TOP LEVEL CELL: Two_bit_adder2{sch}
XNAND_2@0 Cin net@49 net@72 Proj2__NAND_2
XNAND_2@1 A B net@76 Proj2__NAND_2
XNAND_2@2 net@72 net@76 Cout Proj2__NAND_2
XXOR_2@1 A B net@49 Proj2__XOR_2
XXOR_2@2 Cin net@49 Sum Proj2__XOR_2

* Spice Code nodes in cell cell 'Two_bit_adder2{sch}'
VDD VDD 0 DC 3.3
VGND GND 0 DC 0
vin A 0 PULSE(5 0 0 1n 1n 2u 4u)
vin2 B 0 PULSE(5 0 0 1n 1n 1u 2u )
vin3 Cin 0 PULSE(5 0 0 1n 1n 4u 8u)
cload out 0 250fF
.tran 0 10u
.include C:\Electric\C5_models.txt
.END

*** SPICE deck for cell HW3_3{sch} from library project_1_delmaybe
*** Created on Wed Mar 04, 2020 23:22:33
*** Last revised on Wed Mar 04, 2020 23:23:21
*** Written on Wed Mar 04, 2020 23:26:35 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: HW3_3{sch}
Mnmos@0 out A net@38 gnd NMOS L=0.35U W=1.75U
Mnmos@1 net@38 net@2 gnd gnd NMOS L=0.35U W=1.75U
Mnmos@2 out net@5 net@44 gnd NMOS L=0.35U W=1.75U
Mnmos@3 net@44 D gnd gnd NMOS L=0.35U W=1.75U
Mnmos@4 net@2 B gnd gnd NMOS L=0.35U W=1.75U
Mnmos@5 net@5 C gnd gnd NMOS L=0.35U W=1.75U
Mpmos@0 net@24 A vdd vdd PMOS L=0.35U W=1.75U
Mpmos@1 net@24 net@2 vdd vdd PMOS L=0.35U W=1.75U
Mpmos@2 out net@5 net@24 vdd PMOS L=0.35U W=1.75U
Mpmos@3 out D net@24 vdd PMOS L=0.35U W=1.75U
Mpmos@4 net@2 B vdd vdd PMOS L=0.35U W=1.75U
Mpmos@5 net@5 C vdd vdd PMOS L=0.35U W=1.75U

* Spice Code nodes in cell cell 'HW3_3{sch}'
VDD VDD 0 DC 3.3
VGND GND 0 DC 0
vin A 0 PULSE(3.3 0 0 5ns 10ns 100ns 200ns)
vin2 B 0 PULSE(3.3 0 0 5ns 10ns 200ns 400ns)
vin3 C 0 PULSE(3.3 0 0 5ns 10ns 400ns 800ns)
vin4 D 0 PULSE(3.3 0 0 5ns 10ns 800ns 1600ns)
cload out 0 250fF
.tran 0 1600ns
.include C:\Electric\C5_models.txt
.END
